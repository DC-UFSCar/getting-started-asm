module hello()
    // uncomment the following line
    initial
    // $display("Hello, Verilog!");
endmodule